module FechaduraTop (
input 	logic clk, rst, sensor_de_contato, botao_interno,
input	logic [3:0] matricial_col,
output	logic [3:0] matricial_lin,
output 	logic [6:0] dispHex0, dispHex1, dispHex2, dispHex3, dispHex4, dispHex5,
output logic tranca, bip );

endmodule;
